`ifndef AMULET_STATES
`define AMULET_STATES

package amulet_states;
	typedef enum logic [1:0] {A0, A1} amulet_state;
endpackage

`endif