package states;
	typedef enum logic [13:0] {
		FETCH  	= 14'b0_1_0_0_1_10_10_00_0_00,
		DECODE 	= 14'b0_0_0_0_0_00_01_01_0_00,
		MEMADR 	= 14'b0_0_0_0_0_00_01_10_0_00,
		EXECUTER = 14'b0_0_0_0_0_00_00_10_0_10,
		EXECUTEL = 14'b0_0_0_0_0_00_01_10_0_10,
		JAL 		= 14'b0_1_0_0_0_00_10_01_0_00,
		BEQ		= 14'b1_0_0_0_0_00_00_10_0_01,
		MEMREAD  = 14'b0_0_0_0_0_00_00_00_1_00,
		MEMWRITE = 14'b0_0_0_1_0_00_00_00_1_00,
		ALUWB		= 14'b0_0_1_0_0_00_00_00_0_00,
		MEMWB		= 14'b0_0_1_0_0_01_00_00_0_00,
		UNKNOWN  = 14'bx_x_x_x_x_xx_xx_xx_x_xx
	} state;
endpackage