`ifndef GOLD_STATES
`define GOLD_STATES

package gold_states;
	typedef enum logic [1:0] {G0, G1} gold_state;
endpackage

`endif