`ifndef SHIELD_STATES
`define SHIELD_STATES

package shield_states;
	typedef enum logic [1:0] {SH0, SH1} shield_state;
endpackage

`endif