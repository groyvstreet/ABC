`ifndef SWORD_STATES
`define SWORD_STATES

package sword_states;
	typedef enum logic [1:0] {SW0, SW1} sword_state;
endpackage

`endif